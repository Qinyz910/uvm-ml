package mem_env_pkg;
  
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  import mem_agent_pkg::*;
  import mem_sequences_pkg::*;
  
  `include "mem_scoreboard.svh"
  `include "mem_env.svh"

endpackage
