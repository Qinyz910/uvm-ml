package mem_agent_pkg;
  
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  import mem_sequences_pkg::*;
  
  `include "mem_config.svh"
  `include "mem_sequencer.svh"
  `include "mem_driver.svh"
  `include "mem_monitor.svh"
  `include "mem_coverage.svh"
  `include "mem_agent.svh"

endpackage
